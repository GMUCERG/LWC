../../../../LWC_rtl/LWC.vhd