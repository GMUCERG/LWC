../../../LWCsrc/LWC.vhd