../../../LWCsrc/PostProcessor.vhd