../../../../LWCsrc/PreProcessor.vhd