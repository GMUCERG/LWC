../../../LWCsrc/NIST_LWAPI_pkg.vhd