../../../LWCsrc/PreProcessor.vhd