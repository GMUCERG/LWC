../../../../LWC_rtl/StepDownCountLd.vhd