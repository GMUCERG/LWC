../../LWC_tb/LWC_TB.vhd