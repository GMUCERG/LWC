../../../../LWCsrc/fwft_fifo_tb.vhd