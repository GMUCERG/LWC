../../../LWC_rtl/PISO.vhd