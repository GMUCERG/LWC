../../../../LWC_rtl/LWC_wrapper.vhd