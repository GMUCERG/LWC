../../../../LWCsrc/StepDownCountLd.vhd