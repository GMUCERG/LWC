../../../LWC_rtl/SIPO.vhd