../../../LWC_rtl/LWC_pkg.vhd