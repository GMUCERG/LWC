../../../LWCsrc/key_piso.vhd