../../../../LWC_rtl/data_piso.vhd