../../../LWCsrc/data_sipo.vhd