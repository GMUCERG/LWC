../../../../LWC_rtl/fwft_fifo_tb.vhd