../../../LWCsrc/LWC_TB.vhd