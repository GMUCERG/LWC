../../LWC_tb/fwft_fifo_tb.vhd