../../../LWCsrc/StepDownCountLd.vhd