../../../../LWC_rtl/elastic_reg_fifo.vhd