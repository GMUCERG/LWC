../../../LWC_rtl/fifo.vhd