../../LWC_tb/LWC_TB_pkg.vhd