../../../../LWCsrc/LWC.vhd