../../LWC_tb/LWC_TB_compatibility_pkg.vhd