../v1/SPDRam.vhd