../../LWCsrc/lwc_std_logic_1164_additions.vhd