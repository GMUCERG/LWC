../../../LWCsrc/fwft_fifo.vhd