../../../../LWCsrc/PostProcessor.vhd