../../../LWCsrc/data_piso.vhd